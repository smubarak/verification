module tb;

initial $display("Hello HW!");

endmodule
